`include "pyc_handshake_pkg.sv"
`include "pyc_stream_if.sv"
`include "pyc_mem_if.sv"
`include "pyc_add.sv"
`include "pyc_mux.sv"
`include "pyc_and.sv"
`include "pyc_or.sv"
`include "pyc_xor.sv"
`include "pyc_not.sv"
`include "pyc_reg.sv"
`include "pyc_fifo.sv"

`include "pyc_byte_mem.sv"

`include "pyc_queue.sv"
`include "pyc_picker_onehot.sv"
`include "pyc_rr_arb.sv"
`include "pyc_sram.sv"

module linx_cpu_pyc (
  input logic clk,
  input logic rst,
  input logic [63:0] boot_pc,
  input logic [63:0] boot_sp,
  output logic halted,
  output logic [63:0] pc,
  output logic [2:0] stage,
  output logic [63:0] cycles,
  output logic [63:0] a0,
  output logic [63:0] a1,
  output logic [63:0] ra,
  output logic [63:0] sp,
  output logic [1:0] br_kind,
  output logic [63:0] if_window,
  output logic [5:0] wb_op,
  output logic [5:0] wb_regdst,
  output logic [63:0] wb_value,
  output logic commit_cond,
  output logic [63:0] commit_tgt
);

logic [2:0] v1;
logic [1:0] v2;
logic [1:0] v3;
logic [1:0] v4;
logic [63:0] v5;
logic [5:0] v6;
logic [5:0] v7;
logic [5:0] v8;
logic [5:0] v9;
logic [5:0] v10;
logic [2:0] v11;
logic [5:0] v12;
logic [47:0] v13;
logic [47:0] v14;
logic [5:0] v15;
logic [31:0] v16;
logic [31:0] v17;
logic [5:0] v18;
logic [31:0] v19;
logic [31:0] v20;
logic [31:0] v21;
logic [31:0] v22;
logic [5:0] v23;
logic [31:0] v24;
logic [31:0] v25;
logic [5:0] v26;
logic [31:0] v27;
logic [5:0] v28;
logic [31:0] v29;
logic [5:0] v30;
logic [31:0] v31;
logic [5:0] v32;
logic [31:0] v33;
logic [5:0] v34;
logic [31:0] v35;
logic [31:0] v36;
logic [5:0] v37;
logic [31:0] v38;
logic [5:0] v39;
logic [31:0] v40;
logic [5:0] v41;
logic [31:0] v42;
logic [5:0] v43;
logic [31:0] v44;
logic [5:0] v45;
logic [31:0] v46;
logic [31:0] v47;
logic [5:0] v48;
logic [15:0] v49;
logic [5:0] v50;
logic [15:0] v51;
logic [15:0] v52;
logic [5:0] v53;
logic [15:0] v54;
logic [15:0] v55;
logic [15:0] v56;
logic [5:0] v57;
logic [15:0] v58;
logic [5:0] v59;
logic [15:0] v60;
logic [5:0] v61;
logic [15:0] v62;
logic [5:0] v63;
logic [5:0] v64;
logic [15:0] v65;
logic [5:0] v66;
logic [5:0] v67;
logic [15:0] v68;
logic [15:0] v69;
logic [5:0] v70;
logic [15:0] v71;
logic [15:0] v72;
logic [3:0] v73;
logic [7:0] v74;
logic [7:0] v75;
logic [5:0] v76;
logic [2:0] v77;
logic [2:0] v78;
logic [2:0] v79;
logic [2:0] v80;
logic [5:0] v81;
logic [1:0] v82;
logic v83;
logic v84;
logic [2:0] v85;
logic [5:0] v86;
logic [7:0] v87;
logic [63:0] v88;
logic [63:0] v89;
logic [2:0] v90;
logic [1:0] v91;
logic [1:0] v92;
logic [1:0] v93;
logic [63:0] v94;
logic [5:0] v95;
logic [5:0] v96;
logic [5:0] v97;
logic [5:0] v98;
logic [5:0] v99;
logic [2:0] v100;
logic [5:0] v101;
logic [47:0] v102;
logic [47:0] v103;
logic [5:0] v104;
logic [31:0] v105;
logic [31:0] v106;
logic [5:0] v107;
logic [31:0] v108;
logic [31:0] v109;
logic [31:0] v110;
logic [31:0] v111;
logic [5:0] v112;
logic [31:0] v113;
logic [31:0] v114;
logic [5:0] v115;
logic [31:0] v116;
logic [5:0] v117;
logic [31:0] v118;
logic [5:0] v119;
logic [31:0] v120;
logic [5:0] v121;
logic [31:0] v122;
logic [5:0] v123;
logic [31:0] v124;
logic [31:0] v125;
logic [5:0] v126;
logic [31:0] v127;
logic [5:0] v128;
logic [31:0] v129;
logic [5:0] v130;
logic [31:0] v131;
logic [5:0] v132;
logic [31:0] v133;
logic [5:0] v134;
logic [31:0] v135;
logic [31:0] v136;
logic [5:0] v137;
logic [15:0] v138;
logic [5:0] v139;
logic [15:0] v140;
logic [15:0] v141;
logic [5:0] v142;
logic [15:0] v143;
logic [15:0] v144;
logic [15:0] v145;
logic [5:0] v146;
logic [15:0] v147;
logic [5:0] v148;
logic [15:0] v149;
logic [5:0] v150;
logic [15:0] v151;
logic [5:0] v152;
logic [5:0] v153;
logic [15:0] v154;
logic [5:0] v155;
logic [5:0] v156;
logic [15:0] v157;
logic [15:0] v158;
logic [5:0] v159;
logic [15:0] v160;
logic [15:0] v161;
logic [3:0] v162;
logic [7:0] v163;
logic [7:0] v164;
logic [5:0] v165;
logic [2:0] v166;
logic [2:0] v167;
logic [2:0] v168;
logic [2:0] v169;
logic [5:0] v170;
logic [1:0] v171;
logic v172;
logic v173;
logic [2:0] v174;
logic [5:0] v175;
logic [7:0] v176;
logic [63:0] v177;
logic [63:0] v178;
logic [2:0] v179;
logic [2:0] v180;
logic [63:0] v181;
logic [63:0] v182;
logic [1:0] v183;
logic [1:0] v184;
logic [63:0] v185;
logic [63:0] v186;
logic [63:0] v187;
logic [63:0] v188;
logic v189;
logic v190;
logic [63:0] v191;
logic [63:0] v192;
logic [63:0] v193;
logic [63:0] v194;
logic v195;
logic v196;
logic [63:0] v197;
logic [63:0] v198;
logic [5:0] v199;
logic [5:0] v200;
logic [2:0] v201;
logic [2:0] v202;
logic [5:0] v203;
logic [5:0] v204;
logic [5:0] v205;
logic [5:0] v206;
logic [5:0] v207;
logic [5:0] v208;
logic [5:0] v209;
logic [5:0] v210;
logic [63:0] v211;
logic [63:0] v212;
logic [63:0] v213;
logic [63:0] v214;
logic [63:0] v215;
logic [63:0] v216;
logic [63:0] v217;
logic [63:0] v218;
logic [5:0] v219;
logic [5:0] v220;
logic [2:0] v221;
logic [2:0] v222;
logic [5:0] v223;
logic [5:0] v224;
logic [63:0] v225;
logic [63:0] v226;
logic v227;
logic v228;
logic v229;
logic v230;
logic [2:0] v231;
logic [2:0] v232;
logic [63:0] v233;
logic [63:0] v234;
logic [63:0] v235;
logic [63:0] v236;
logic [5:0] v237;
logic [5:0] v238;
logic [2:0] v239;
logic [2:0] v240;
logic [5:0] v241;
logic [5:0] v242;
logic [63:0] v243;
logic [63:0] v244;
logic [63:0] v245;
logic [63:0] v246;
logic [63:0] v247;
logic [63:0] v248;
logic [63:0] v249;
logic [63:0] v250;
logic [63:0] v251;
logic [63:0] v252;
logic [63:0] v253;
logic [63:0] v254;
logic [63:0] v255;
logic [63:0] v256;
logic [63:0] v257;
logic [63:0] v258;
logic [63:0] v259;
logic [63:0] v260;
logic [63:0] v261;
logic [63:0] v262;
logic [63:0] v263;
logic [63:0] v264;
logic [63:0] v265;
logic [63:0] v266;
logic [63:0] v267;
logic [63:0] v268;
logic [63:0] v269;
logic [63:0] v270;
logic [63:0] v271;
logic [63:0] v272;
logic [63:0] v273;
logic [63:0] v274;
logic [63:0] v275;
logic [63:0] v276;
logic [63:0] v277;
logic [63:0] v278;
logic [63:0] v279;
logic [63:0] v280;
logic [63:0] v281;
logic [63:0] v282;
logic [63:0] v283;
logic [63:0] v284;
logic [63:0] v285;
logic [63:0] v286;
logic [63:0] v287;
logic [63:0] v288;
logic [63:0] v289;
logic [63:0] v290;
logic [63:0] v291;
logic [63:0] v292;
logic [63:0] v293;
logic [63:0] v294;
logic [63:0] v295;
logic [63:0] v296;
logic [63:0] v297;
logic [63:0] v298;
logic [63:0] v299;
logic [63:0] v300;
logic [63:0] v301;
logic [63:0] v302;
logic [63:0] v303;
logic [63:0] v304;
logic [63:0] v305;
logic [63:0] v306;
logic [63:0] v307;
logic [63:0] v308;
logic v309;
logic v310;
logic v311;
logic v312;
logic v313;
logic v314;
logic v315;
logic v316;
logic v317;
logic v318;
logic v319;
logic v320;
logic v321;
logic v322;
logic v323;
logic v324;
logic v325;
logic v326;
logic v327;
logic [63:0] v328;
logic [63:0] v329;
logic v330;
logic v331;
logic [7:0] v332;
logic v333;
logic [7:0] v334;
logic v335;
logic v336;
logic v337;
logic v338;
logic v339;
logic v340;
logic v341;
logic v342;
logic v343;
logic v344;
logic v345;
logic v346;
logic [63:0] v347;
logic v348;
logic [7:0] v349;
logic [63:0] v350;
logic [63:0] v351;
logic [15:0] v352;
logic [31:0] v353;
logic [47:0] v354;
logic [3:0] v355;
logic v356;
logic v357;
logic v358;
logic v359;
logic v360;
logic v361;
logic [4:0] v362;
logic [5:0] v363;
logic [4:0] v364;
logic [5:0] v365;
logic [4:0] v366;
logic [5:0] v367;
logic [4:0] v368;
logic [5:0] v369;
logic [11:0] v370;
logic [63:0] v371;
logic [63:0] v372;
logic [19:0] v373;
logic [63:0] v374;
logic [6:0] v375;
logic [11:0] v376;
logic [11:0] v377;
logic [11:0] v378;
logic [11:0] v379;
logic [63:0] v380;
logic [16:0] v381;
logic [63:0] v382;
logic [15:0] v383;
logic [31:0] v384;
logic [11:0] v385;
logic [19:0] v386;
logic [31:0] v387;
logic [31:0] v388;
logic [31:0] v389;
logic [31:0] v390;
logic [63:0] v391;
logic [4:0] v392;
logic [5:0] v393;
logic [4:0] v394;
logic [5:0] v395;
logic [4:0] v396;
logic [5:0] v397;
logic [63:0] v398;
logic [63:0] v399;
logic [11:0] v400;
logic [63:0] v401;
logic [63:0] v402;
logic [2:0] v403;
logic [63:0] v404;
logic [15:0] v405;
logic v406;
logic v407;
logic [5:0] v408;
logic [2:0] v409;
logic [5:0] v410;
logic [5:0] v411;
logic [63:0] v412;
logic [15:0] v413;
logic v414;
logic v415;
logic [63:0] v416;
logic [5:0] v417;
logic [2:0] v418;
logic [5:0] v419;
logic [5:0] v420;
logic [63:0] v421;
logic v422;
logic v423;
logic [5:0] v424;
logic [2:0] v425;
logic [5:0] v426;
logic [5:0] v427;
logic [5:0] v428;
logic [5:0] v429;
logic [63:0] v430;
logic v431;
logic v432;
logic [5:0] v433;
logic [2:0] v434;
logic [5:0] v435;
logic [5:0] v436;
logic [5:0] v437;
logic [5:0] v438;
logic [63:0] v439;
logic v440;
logic v441;
logic [5:0] v442;
logic [2:0] v443;
logic [5:0] v444;
logic [5:0] v445;
logic [5:0] v446;
logic [5:0] v447;
logic [63:0] v448;
logic v449;
logic v450;
logic [5:0] v451;
logic [2:0] v452;
logic [5:0] v453;
logic [5:0] v454;
logic [5:0] v455;
logic [5:0] v456;
logic [63:0] v457;
logic v458;
logic v459;
logic [5:0] v460;
logic [2:0] v461;
logic [5:0] v462;
logic [5:0] v463;
logic [5:0] v464;
logic [5:0] v465;
logic [63:0] v466;
logic [15:0] v467;
logic v468;
logic v469;
logic [63:0] v470;
logic [5:0] v471;
logic [2:0] v472;
logic [5:0] v473;
logic [5:0] v474;
logic [5:0] v475;
logic [5:0] v476;
logic [63:0] v477;
logic [15:0] v478;
logic v479;
logic v480;
logic [5:0] v481;
logic [2:0] v482;
logic [5:0] v483;
logic [5:0] v484;
logic [5:0] v485;
logic [5:0] v486;
logic [63:0] v487;
logic [15:0] v488;
logic v489;
logic v490;
logic [5:0] v491;
logic [2:0] v492;
logic [5:0] v493;
logic [5:0] v494;
logic [5:0] v495;
logic [5:0] v496;
logic [63:0] v497;
logic [31:0] v498;
logic v499;
logic v500;
logic [5:0] v501;
logic [2:0] v502;
logic [5:0] v503;
logic [5:0] v504;
logic [5:0] v505;
logic [5:0] v506;
logic [63:0] v507;
logic v508;
logic v509;
logic [5:0] v510;
logic [2:0] v511;
logic [5:0] v512;
logic [5:0] v513;
logic [5:0] v514;
logic [5:0] v515;
logic [63:0] v516;
logic v517;
logic v518;
logic [5:0] v519;
logic [2:0] v520;
logic [5:0] v521;
logic [5:0] v522;
logic [5:0] v523;
logic [5:0] v524;
logic [63:0] v525;
logic v526;
logic v527;
logic [5:0] v528;
logic [2:0] v529;
logic [5:0] v530;
logic [5:0] v531;
logic [5:0] v532;
logic [5:0] v533;
logic [63:0] v534;
logic v535;
logic v536;
logic [5:0] v537;
logic [2:0] v538;
logic [5:0] v539;
logic [5:0] v540;
logic [5:0] v541;
logic [5:0] v542;
logic [63:0] v543;
logic v544;
logic v545;
logic [5:0] v546;
logic [2:0] v547;
logic [5:0] v548;
logic [5:0] v549;
logic [5:0] v550;
logic [5:0] v551;
logic [63:0] v552;
logic v553;
logic v554;
logic [5:0] v555;
logic [2:0] v556;
logic [5:0] v557;
logic [5:0] v558;
logic [5:0] v559;
logic [5:0] v560;
logic [63:0] v561;
logic v562;
logic v563;
logic [5:0] v564;
logic [2:0] v565;
logic [5:0] v566;
logic [5:0] v567;
logic [5:0] v568;
logic [5:0] v569;
logic [63:0] v570;
logic v571;
logic v572;
logic [5:0] v573;
logic [2:0] v574;
logic [5:0] v575;
logic [5:0] v576;
logic [5:0] v577;
logic [5:0] v578;
logic [63:0] v579;
logic v580;
logic v581;
logic [5:0] v582;
logic [2:0] v583;
logic [5:0] v584;
logic [5:0] v585;
logic [5:0] v586;
logic [5:0] v587;
logic [63:0] v588;
logic v589;
logic v590;
logic [5:0] v591;
logic [2:0] v592;
logic [5:0] v593;
logic [5:0] v594;
logic [5:0] v595;
logic [5:0] v596;
logic [63:0] v597;
logic [31:0] v598;
logic v599;
logic v600;
logic [5:0] v601;
logic [2:0] v602;
logic [5:0] v603;
logic [5:0] v604;
logic [5:0] v605;
logic [5:0] v606;
logic [63:0] v607;
logic [31:0] v608;
logic v609;
logic v610;
logic [5:0] v611;
logic [2:0] v612;
logic [5:0] v613;
logic [5:0] v614;
logic [5:0] v615;
logic [5:0] v616;
logic [63:0] v617;
logic [31:0] v618;
logic v619;
logic v620;
logic [63:0] v621;
logic [5:0] v622;
logic [2:0] v623;
logic [5:0] v624;
logic [5:0] v625;
logic [5:0] v626;
logic [5:0] v627;
logic [63:0] v628;
logic [31:0] v629;
logic v630;
logic v631;
logic [63:0] v632;
logic [5:0] v633;
logic [2:0] v634;
logic [5:0] v635;
logic [5:0] v636;
logic [5:0] v637;
logic [5:0] v638;
logic [63:0] v639;
logic [47:0] v640;
logic v641;
logic v642;
logic [5:0] v643;
logic [2:0] v644;
logic [5:0] v645;
logic [5:0] v646;
logic [5:0] v647;
logic [5:0] v648;
logic [63:0] v649;
logic [5:0] v650;
logic [2:0] v651;
logic [5:0] v652;
logic [5:0] v653;
logic [5:0] v654;
logic [5:0] v655;
logic [63:0] v656;
logic [5:0] v657;
logic [2:0] v658;
logic [5:0] v659;
logic [5:0] v660;
logic [5:0] v661;
logic [5:0] v662;
logic [63:0] v663;
logic v664;
logic [63:0] v665;
logic v666;
logic [63:0] v667;
logic v668;
logic [63:0] v669;
logic v670;
logic [63:0] v671;
logic v672;
logic [63:0] v673;
logic v674;
logic [63:0] v675;
logic v676;
logic [63:0] v677;
logic v678;
logic [63:0] v679;
logic v680;
logic [63:0] v681;
logic v682;
logic [63:0] v683;
logic v684;
logic [63:0] v685;
logic v686;
logic [63:0] v687;
logic v688;
logic [63:0] v689;
logic v690;
logic [63:0] v691;
logic v692;
logic [63:0] v693;
logic v694;
logic [63:0] v695;
logic v696;
logic [63:0] v697;
logic v698;
logic [63:0] v699;
logic v700;
logic [63:0] v701;
logic v702;
logic [63:0] v703;
logic v704;
logic [63:0] v705;
logic v706;
logic [63:0] v707;
logic v708;
logic [63:0] v709;
logic v710;
logic [63:0] v711;
logic v712;
logic [63:0] v713;
logic v714;
logic [63:0] v715;
logic v716;
logic [63:0] v717;
logic v718;
logic [63:0] v719;
logic v720;
logic [63:0] v721;
logic v722;
logic [63:0] v723;
logic v724;
logic [63:0] v725;
logic v726;
logic [63:0] v727;
logic v728;
logic [63:0] v729;
logic v730;
logic [63:0] v731;
logic v732;
logic [63:0] v733;
logic v734;
logic [63:0] v735;
logic v736;
logic [63:0] v737;
logic v738;
logic [63:0] v739;
logic v740;
logic [63:0] v741;
logic v742;
logic [63:0] v743;
logic v744;
logic [63:0] v745;
logic v746;
logic [63:0] v747;
logic v748;
logic [63:0] v749;
logic v750;
logic [63:0] v751;
logic v752;
logic [63:0] v753;
logic v754;
logic [63:0] v755;
logic v756;
logic [63:0] v757;
logic v758;
logic [63:0] v759;
logic v760;
logic [63:0] v761;
logic v762;
logic [63:0] v763;
logic v764;
logic [63:0] v765;
logic v766;
logic [63:0] v767;
logic v768;
logic [63:0] v769;
logic v770;
logic [63:0] v771;
logic v772;
logic [63:0] v773;
logic v774;
logic [63:0] v775;
logic v776;
logic [63:0] v777;
logic v778;
logic [63:0] v779;
logic v780;
logic [63:0] v781;
logic v782;
logic [63:0] v783;
logic v784;
logic [63:0] v785;
logic v786;
logic [63:0] v787;
logic v788;
logic [63:0] v789;
logic v790;
logic [63:0] v791;
logic v792;
logic [63:0] v793;
logic v794;
logic [63:0] v795;
logic v796;
logic [63:0] v797;
logic v798;
logic [63:0] v799;
logic v800;
logic [63:0] v801;
logic v802;
logic [63:0] v803;
logic v804;
logic [63:0] v805;
logic v806;
logic [63:0] v807;
logic v808;
logic [63:0] v809;
logic v810;
logic [63:0] v811;
logic v812;
logic [63:0] v813;
logic v814;
logic [63:0] v815;
logic v816;
logic [63:0] v817;
logic v818;
logic [63:0] v819;
logic v820;
logic [63:0] v821;
logic v822;
logic [63:0] v823;
logic v824;
logic [63:0] v825;
logic v826;
logic [63:0] v827;
logic v828;
logic [63:0] v829;
logic v830;
logic [63:0] v831;
logic v832;
logic [63:0] v833;
logic v834;
logic [63:0] v835;
logic v836;
logic [63:0] v837;
logic v838;
logic [63:0] v839;
logic v840;
logic [63:0] v841;
logic v842;
logic [63:0] v843;
logic v844;
logic [63:0] v845;
logic v846;
logic [63:0] v847;
logic v848;
logic [63:0] v849;
logic v850;
logic [63:0] v851;
logic v852;
logic [63:0] v853;
logic v854;
logic [63:0] v855;
logic [63:0] v856;
logic [63:0] v857;
logic [63:0] v858;
logic [63:0] v859;
logic [63:0] v860;
logic [63:0] v861;
logic v862;
logic v863;
logic v864;
logic v865;
logic v866;
logic v867;
logic v868;
logic v869;
logic v870;
logic v871;
logic v872;
logic v873;
logic v874;
logic v875;
logic v876;
logic v877;
logic v878;
logic v879;
logic v880;
logic v881;
logic v882;
logic v883;
logic v884;
logic v885;
logic [63:0] v886;
logic v887;
logic v888;
logic [63:0] v889;
logic v890;
logic [2:0] v891;
logic [63:0] v892;
logic [63:0] v893;
logic v894;
logic [2:0] v895;
logic [63:0] v896;
logic [63:0] v897;
logic v898;
logic [2:0] v899;
logic [63:0] v900;
logic [63:0] v901;
logic [63:0] v902;
logic v903;
logic [2:0] v904;
logic [63:0] v905;
logic v906;
logic [63:0] v907;
logic [63:0] v908;
logic v909;
logic [2:0] v910;
logic [63:0] v911;
logic [63:0] v912;
logic v913;
logic [2:0] v914;
logic [63:0] v915;
logic [63:0] v916;
logic [63:0] v917;
logic [63:0] v918;
logic v919;
logic [2:0] v920;
logic [63:0] v921;
logic [63:0] v922;
logic [63:0] v923;
logic v924;
logic [2:0] v925;
logic [63:0] v926;
logic [63:0] v927;
logic [63:0] v928;
logic [63:0] v929;
logic [63:0] v930;
logic v931;
logic [2:0] v932;
logic [63:0] v933;
logic [31:0] v934;
logic [31:0] v935;
logic [31:0] v936;
logic [63:0] v937;
logic [63:0] v938;
logic v939;
logic [2:0] v940;
logic [63:0] v941;
logic [31:0] v942;
logic [31:0] v943;
logic [63:0] v944;
logic [31:0] v945;
logic [63:0] v946;
logic [31:0] v947;
logic [63:0] v948;
logic [31:0] v949;
logic [63:0] v950;
logic [63:0] v951;
logic v952;
logic [2:0] v953;
logic [63:0] v954;
logic [63:0] v955;
logic v956;
logic [2:0] v957;
logic [63:0] v958;
logic [63:0] v959;
logic v960;
logic [2:0] v961;
logic [63:0] v962;
logic [63:0] v963;
logic v964;
logic [2:0] v965;
logic [63:0] v966;
logic [63:0] v967;
logic v968;
logic [2:0] v969;
logic [63:0] v970;
logic [63:0] v971;
logic v972;
logic [2:0] v973;
logic [63:0] v974;
logic v975;
logic v976;
logic [63:0] v977;
logic [63:0] v978;
logic v979;
logic [2:0] v980;
logic [63:0] v981;
logic v982;
logic [63:0] v983;
logic [63:0] v984;
logic v985;
logic v986;
logic [2:0] v987;
logic [63:0] v988;
logic [63:0] v989;
logic [63:0] v990;
logic [63:0] v991;
logic [63:0] v992;
logic v993;
logic [63:0] v994;
logic v995;
logic v996;
logic [2:0] v997;
logic [63:0] v998;
logic [63:0] v999;
logic [63:0] v1000;
logic [63:0] v1001;
logic [63:0] v1002;
logic v1003;
logic v1004;
logic [2:0] v1005;
logic [63:0] v1006;
logic [63:0] v1007;
logic [5:0] v1008;
logic [63:0] v1009;
logic v1010;
logic v1011;
logic [2:0] v1012;
logic [63:0] v1013;
logic [63:0] v1014;
logic [5:0] v1015;
logic [2:0] v1016;
logic [5:0] v1017;
logic [63:0] v1018;
logic v1019;
logic v1020;
logic [2:0] v1021;
logic [63:0] v1022;
logic [63:0] v1023;
logic [31:0] v1024;
logic [63:0] v1025;
logic [63:0] v1026;
logic [63:0] v1027;
logic [5:0] v1028;
logic [63:0] v1029;
logic [5:0] v1030;
logic [2:0] v1031;
logic [5:0] v1032;
logic [63:0] v1033;
logic v1034;
logic v1035;
logic v1036;
logic v1037;
logic v1038;
logic v1039;
logic v1040;
logic v1041;
logic v1042;
logic v1043;
logic v1044;
logic [63:0] v1045;
logic [63:0] v1046;
logic v1047;
logic v1048;
logic v1049;
logic [63:0] v1050;
logic [63:0] v1051;
logic [63:0] v1052;
logic [63:0] v1053;
logic [63:0] v1054;
logic v1055;
logic v1056;
logic v1057;
logic v1058;
logic v1059;
logic v1060;
logic v1061;
logic [63:0] v1062;
logic [2:0] v1063;
logic [2:0] v1064;
logic [2:0] v1065;
logic [2:0] v1066;
logic [2:0] v1067;
logic [2:0] v1068;
logic [2:0] v1069;
logic [63:0] v1070;
logic v1071;
logic v1072;
logic v1073;
logic v1074;
logic [63:0] v1075;
logic v1076;
logic v1077;
logic v1078;
logic v1079;
logic [63:0] v1080;
logic v1081;
logic v1082;
logic [63:0] v1083;
logic v1084;
logic [1:0] v1085;
logic [63:0] v1086;
logic [63:0] v1087;
logic v1088;
logic v1089;
logic v1090;
logic v1091;
logic [1:0] v1092;
logic [63:0] v1093;
logic [63:0] v1094;
logic v1095;
logic [1:0] v1096;
logic [63:0] v1097;
logic [63:0] v1098;
logic [2:0] v1099;
logic v1100;
logic [1:0] v1101;
logic v1102;
logic [1:0] v1103;
logic [63:0] v1104;
logic [63:0] v1105;
logic v1106;
logic [1:0] v1107;
logic [63:0] v1108;
logic [63:0] v1109;
logic v1110;
logic [1:0] v1111;
logic [63:0] v1112;
logic [63:0] v1113;
logic v1114;
logic v1115;
logic v1116;
logic v1117;
logic v1118;
logic v1119;
logic v1120;
logic v1121;
logic v1122;
logic v1123;
logic v1124;
logic v1125;
logic v1126;
logic v1127;
logic v1128;
logic v1129;
logic v1130;
logic v1131;
logic v1132;
logic v1133;
logic [63:0] v1134;
logic [63:0] v1135;
logic v1136;
logic v1137;
logic [63:0] v1138;
logic [63:0] v1139;
logic v1140;
logic v1141;
logic [63:0] v1142;
logic [63:0] v1143;
logic v1144;
logic v1145;
logic [63:0] v1146;
logic [63:0] v1147;
logic v1148;
logic v1149;
logic [63:0] v1150;
logic [63:0] v1151;
logic v1152;
logic v1153;
logic [63:0] v1154;
logic [63:0] v1155;
logic v1156;
logic v1157;
logic [63:0] v1158;
logic [63:0] v1159;
logic v1160;
logic v1161;
logic [63:0] v1162;
logic [63:0] v1163;
logic v1164;
logic v1165;
logic [63:0] v1166;
logic [63:0] v1167;
logic v1168;
logic v1169;
logic [63:0] v1170;
logic [63:0] v1171;
logic v1172;
logic v1173;
logic [63:0] v1174;
logic [63:0] v1175;
logic v1176;
logic v1177;
logic [63:0] v1178;
logic [63:0] v1179;
logic v1180;
logic v1181;
logic [63:0] v1182;
logic [63:0] v1183;
logic v1184;
logic v1185;
logic [63:0] v1186;
logic [63:0] v1187;
logic v1188;
logic v1189;
logic [63:0] v1190;
logic [63:0] v1191;
logic v1192;
logic v1193;
logic [63:0] v1194;
logic [63:0] v1195;
logic v1196;
logic v1197;
logic [63:0] v1198;
logic [63:0] v1199;
logic v1200;
logic v1201;
logic [63:0] v1202;
logic [63:0] v1203;
logic v1204;
logic v1205;
logic [63:0] v1206;
logic [63:0] v1207;
logic v1208;
logic v1209;
logic [63:0] v1210;
logic [63:0] v1211;
logic v1212;
logic v1213;
logic [63:0] v1214;
logic [63:0] v1215;
logic v1216;
logic v1217;
logic [63:0] v1218;
logic [63:0] v1219;
logic v1220;
logic v1221;
logic [63:0] v1222;
logic [63:0] v1223;
logic [63:0] v1224;
logic [63:0] v1225;
logic [63:0] v1226;
logic [63:0] v1227;
logic [63:0] v1228;
logic [63:0] v1229;
logic [63:0] v1230;
logic [63:0] v1231;
logic [63:0] v1232;
logic [63:0] v1233;
logic [63:0] v1234;
logic [63:0] v1235;
logic [63:0] v1236;
logic [63:0] v1237;
logic [63:0] v1238;
logic [63:0] v1239;
logic [63:0] v1240;
logic [63:0] v1241;
logic [63:0] v1242;
logic [63:0] v1243;
logic [63:0] v1244;
logic [63:0] v1245;
logic [63:0] v1246;
logic [63:0] v1247;

assign v1 = 3'd7;
assign v2 = 2'd3;
assign v3 = 2'd2;
assign v4 = 2'd1;
assign v5 = 64'd18446744073709547520;
assign v6 = 6'd31;
assign v7 = 6'd30;
assign v8 = 6'd29;
assign v9 = 6'd28;
assign v10 = 6'd27;
assign v11 = 3'd6;
assign v12 = 6'd17;
assign v13 = 48'd1507342;
assign v14 = 48'd8323087;
assign v15 = 6'd20;
assign v16 = 32'd16385;
assign v17 = 32'd32767;
assign v18 = 6'd25;
assign v19 = 32'd7;
assign v20 = 32'd127;
assign v21 = 32'd1052715;
assign v22 = 32'd4043309055;
assign v23 = 6'd15;
assign v24 = 32'd69;
assign v25 = 32'd4160778367;
assign v26 = 6'd6;
assign v27 = 32'd4117;
assign v28 = 6'd7;
assign v29 = 32'd21;
assign v30 = 6'd8;
assign v31 = 32'd53;
assign v32 = 6'd9;
assign v33 = 32'd8217;
assign v34 = 6'd26;
assign v35 = 32'd12377;
assign v36 = 32'd8281;
assign v37 = 6'd16;
assign v38 = 32'd119;
assign v39 = 6'd11;
assign v40 = 32'd37;
assign v41 = 6'd12;
assign v42 = 32'd12325;
assign v43 = 6'd13;
assign v44 = 32'd8229;
assign v45 = 6'd14;
assign v46 = 32'd16421;
assign v47 = 32'd28799;
assign v48 = 6'd2;
assign v49 = 16'd65535;
assign v50 = 6'd1;
assign v51 = 16'd0;
assign v52 = 16'd51199;
assign v53 = 6'd19;
assign v54 = 16'd4;
assign v55 = 16'd15;
assign v56 = 16'd28;
assign v57 = 6'd23;
assign v58 = 16'd38;
assign v59 = 6'd3;
assign v60 = 16'd6;
assign v61 = 6'd4;
assign v62 = 16'd10;
assign v63 = 6'd5;
assign v64 = 6'd24;
assign v65 = 16'd42;
assign v66 = 6'd22;
assign v67 = 6'd10;
assign v68 = 16'd20502;
assign v69 = 16'd63551;
assign v70 = 6'd21;
assign v71 = 16'd22;
assign v72 = 16'd63;
assign v73 = 4'd14;
assign v74 = 8'd15;
assign v75 = 8'd255;
assign v76 = 6'd18;
assign v77 = 3'd4;
assign v78 = 3'd3;
assign v79 = 3'd2;
assign v80 = 3'd1;
assign v81 = 6'd63;
assign v82 = 2'd0;
assign v83 = 1'd1;
assign v84 = 1'd0;
assign v85 = 3'd0;
assign v86 = 6'd0;
assign v87 = 8'd0;
assign v88 = 64'd0;
assign v89 = 64'd1;
assign v90 = v1;
assign v91 = v2;
assign v92 = v3;
assign v93 = v4;
assign v94 = v5;
assign v95 = v6;
assign v96 = v7;
assign v97 = v8;
assign v98 = v9;
assign v99 = v10;
assign v100 = v11;
assign v101 = v12;
assign v102 = v13;
assign v103 = v14;
assign v104 = v15;
assign v105 = v16;
assign v106 = v17;
assign v107 = v18;
assign v108 = v19;
assign v109 = v20;
assign v110 = v21;
assign v111 = v22;
assign v112 = v23;
assign v113 = v24;
assign v114 = v25;
assign v115 = v26;
assign v116 = v27;
assign v117 = v28;
assign v118 = v29;
assign v119 = v30;
assign v120 = v31;
assign v121 = v32;
assign v122 = v33;
assign v123 = v34;
assign v124 = v35;
assign v125 = v36;
assign v126 = v37;
assign v127 = v38;
assign v128 = v39;
assign v129 = v40;
assign v130 = v41;
assign v131 = v42;
assign v132 = v43;
assign v133 = v44;
assign v134 = v45;
assign v135 = v46;
assign v136 = v47;
assign v137 = v48;
assign v138 = v49;
assign v139 = v50;
assign v140 = v51;
assign v141 = v52;
assign v142 = v53;
assign v143 = v54;
assign v144 = v55;
assign v145 = v56;
assign v146 = v57;
assign v147 = v58;
assign v148 = v59;
assign v149 = v60;
assign v150 = v61;
assign v151 = v62;
assign v152 = v63;
assign v153 = v64;
assign v154 = v65;
assign v155 = v66;
assign v156 = v67;
assign v157 = v68;
assign v158 = v69;
assign v159 = v70;
assign v160 = v71;
assign v161 = v72;
assign v162 = v73;
assign v163 = v74;
assign v164 = v75;
assign v165 = v76;
assign v166 = v77;
assign v167 = v78;
assign v168 = v79;
assign v169 = v80;
assign v170 = v81;
assign v171 = v82;
assign v172 = v83;
assign v173 = v84;
assign v174 = v85;
assign v175 = v86;
assign v176 = v87;
assign v177 = v88;
assign v178 = v89;
pyc_reg #(.WIDTH(3)) v180_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v179),
  .init(v174),
  .q(v180)
);
pyc_reg #(.WIDTH(64)) v182_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v181),
  .init(boot_pc),
  .q(v182)
);
pyc_reg #(.WIDTH(2)) v184_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v183),
  .init(v171),
  .q(v184)
);
pyc_reg #(.WIDTH(64)) v186_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v185),
  .init(boot_pc),
  .q(v186)
);
pyc_reg #(.WIDTH(64)) v188_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v187),
  .init(v177),
  .q(v188)
);
pyc_reg #(.WIDTH(1)) v190_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v189),
  .init(v173),
  .q(v190)
);
pyc_reg #(.WIDTH(64)) v192_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v191),
  .init(v177),
  .q(v192)
);
pyc_reg #(.WIDTH(64)) v194_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v193),
  .init(v177),
  .q(v194)
);
pyc_reg #(.WIDTH(1)) v196_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v195),
  .init(v173),
  .q(v196)
);
pyc_reg #(.WIDTH(64)) v198_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v197),
  .init(v177),
  .q(v198)
);
pyc_reg #(.WIDTH(6)) v200_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v199),
  .init(v175),
  .q(v200)
);
pyc_reg #(.WIDTH(3)) v202_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v201),
  .init(v174),
  .q(v202)
);
pyc_reg #(.WIDTH(6)) v204_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v203),
  .init(v170),
  .q(v204)
);
pyc_reg #(.WIDTH(6)) v206_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v205),
  .init(v170),
  .q(v206)
);
pyc_reg #(.WIDTH(6)) v208_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v207),
  .init(v170),
  .q(v208)
);
pyc_reg #(.WIDTH(6)) v210_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v209),
  .init(v170),
  .q(v210)
);
pyc_reg #(.WIDTH(64)) v212_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v211),
  .init(v177),
  .q(v212)
);
pyc_reg #(.WIDTH(64)) v214_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v213),
  .init(v177),
  .q(v214)
);
pyc_reg #(.WIDTH(64)) v216_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v215),
  .init(v177),
  .q(v216)
);
pyc_reg #(.WIDTH(64)) v218_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v217),
  .init(v177),
  .q(v218)
);
pyc_reg #(.WIDTH(6)) v220_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v219),
  .init(v175),
  .q(v220)
);
pyc_reg #(.WIDTH(3)) v222_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v221),
  .init(v174),
  .q(v222)
);
pyc_reg #(.WIDTH(6)) v224_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v223),
  .init(v170),
  .q(v224)
);
pyc_reg #(.WIDTH(64)) v226_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v225),
  .init(v177),
  .q(v226)
);
pyc_reg #(.WIDTH(1)) v228_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v227),
  .init(v173),
  .q(v228)
);
pyc_reg #(.WIDTH(1)) v230_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v229),
  .init(v173),
  .q(v230)
);
pyc_reg #(.WIDTH(3)) v232_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v231),
  .init(v174),
  .q(v232)
);
pyc_reg #(.WIDTH(64)) v234_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v233),
  .init(v177),
  .q(v234)
);
pyc_reg #(.WIDTH(64)) v236_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v235),
  .init(v177),
  .q(v236)
);
pyc_reg #(.WIDTH(6)) v238_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v237),
  .init(v175),
  .q(v238)
);
pyc_reg #(.WIDTH(3)) v240_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v239),
  .init(v174),
  .q(v240)
);
pyc_reg #(.WIDTH(6)) v242_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v241),
  .init(v170),
  .q(v242)
);
pyc_reg #(.WIDTH(64)) v244_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v243),
  .init(v177),
  .q(v244)
);
pyc_reg #(.WIDTH(64)) v246_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v245),
  .init(v177),
  .q(v246)
);
pyc_reg #(.WIDTH(64)) v248_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v247),
  .init(boot_sp),
  .q(v248)
);
pyc_reg #(.WIDTH(64)) v250_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v249),
  .init(v177),
  .q(v250)
);
pyc_reg #(.WIDTH(64)) v252_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v251),
  .init(v177),
  .q(v252)
);
pyc_reg #(.WIDTH(64)) v254_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v253),
  .init(v177),
  .q(v254)
);
pyc_reg #(.WIDTH(64)) v256_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v255),
  .init(v177),
  .q(v256)
);
pyc_reg #(.WIDTH(64)) v258_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v257),
  .init(v177),
  .q(v258)
);
pyc_reg #(.WIDTH(64)) v260_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v259),
  .init(v177),
  .q(v260)
);
pyc_reg #(.WIDTH(64)) v262_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v261),
  .init(v177),
  .q(v262)
);
pyc_reg #(.WIDTH(64)) v264_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v263),
  .init(v177),
  .q(v264)
);
pyc_reg #(.WIDTH(64)) v266_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v265),
  .init(v177),
  .q(v266)
);
pyc_reg #(.WIDTH(64)) v268_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v267),
  .init(v177),
  .q(v268)
);
pyc_reg #(.WIDTH(64)) v270_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v269),
  .init(v177),
  .q(v270)
);
pyc_reg #(.WIDTH(64)) v272_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v271),
  .init(v177),
  .q(v272)
);
pyc_reg #(.WIDTH(64)) v274_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v273),
  .init(v177),
  .q(v274)
);
pyc_reg #(.WIDTH(64)) v276_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v275),
  .init(v177),
  .q(v276)
);
pyc_reg #(.WIDTH(64)) v278_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v277),
  .init(v177),
  .q(v278)
);
pyc_reg #(.WIDTH(64)) v280_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v279),
  .init(v177),
  .q(v280)
);
pyc_reg #(.WIDTH(64)) v282_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v281),
  .init(v177),
  .q(v282)
);
pyc_reg #(.WIDTH(64)) v284_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v283),
  .init(v177),
  .q(v284)
);
pyc_reg #(.WIDTH(64)) v286_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v285),
  .init(v177),
  .q(v286)
);
pyc_reg #(.WIDTH(64)) v288_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v287),
  .init(v177),
  .q(v288)
);
pyc_reg #(.WIDTH(64)) v290_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v289),
  .init(v177),
  .q(v290)
);
pyc_reg #(.WIDTH(64)) v292_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v291),
  .init(v177),
  .q(v292)
);
pyc_reg #(.WIDTH(64)) v294_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v293),
  .init(v177),
  .q(v294)
);
pyc_reg #(.WIDTH(64)) v296_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v295),
  .init(v177),
  .q(v296)
);
pyc_reg #(.WIDTH(64)) v298_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v297),
  .init(v177),
  .q(v298)
);
pyc_reg #(.WIDTH(64)) v300_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v299),
  .init(v177),
  .q(v300)
);
pyc_reg #(.WIDTH(64)) v302_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v301),
  .init(v177),
  .q(v302)
);
pyc_reg #(.WIDTH(64)) v304_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v303),
  .init(v177),
  .q(v304)
);
pyc_reg #(.WIDTH(64)) v306_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v305),
  .init(v177),
  .q(v306)
);
pyc_reg #(.WIDTH(64)) v308_inst (
  .clk(clk),
  .rst(rst),
  .en(v172),
  .d(v307),
  .init(v177),
  .q(v308)
);
assign v309 = (v180 == v174);
assign v310 = (v180 == v169);
assign v311 = (v180 == v168);
assign v312 = (v180 == v167);
assign v313 = (v180 == v166);
assign v314 = (~v196);
assign v315 = (v313 & v314);
assign v316 = (v238 == v165);
assign v317 = (v238 == v175);
assign v318 = (v316 | v317);
assign v319 = (v315 & v318);
assign v320 = (v196 | v319);
assign v321 = (~v320);
assign v322 = (v309 & v321);
assign v323 = (v310 & v321);
assign v324 = (v311 & v321);
assign v325 = (v312 & v321);
assign v326 = (v313 & v321);
assign v327 = (v325 & v228);
assign v328 = (v327 ? v234 : v177);
assign v329 = (v322 ? v182 : v328);
assign v330 = (v325 & v230);
assign v331 = (v232 == v174);
assign v332 = (v331 ? v164 : v176);
assign v333 = (v232 == v166);
assign v334 = (v333 ? v163 : v332);
assign v335 = v309;
assign v336 = v310;
assign v337 = v311;
assign v338 = v312;
assign v339 = v313;
assign v340 = v319;
assign v341 = v320;
assign v342 = v322;
assign v343 = v323;
assign v344 = v324;
assign v345 = v325;
assign v346 = v326;
assign v347 = v329;
assign v348 = v330;
assign v349 = v334;
pyc_byte_mem #(.ADDR_WIDTH(64), .DATA_WIDTH(64), .DEPTH(1048576)) mem (
  .clk(clk),
  .rst(rst),
  .raddr(v347),
  .rdata(v350),
  .wvalid(v348),
  .waddr(v234),
  .wdata(v236),
  .wstrb(v349)
);
pyc_mux #(.WIDTH(64)) v351_inst (
  .sel(v342),
  .a(v350),
  .b(v198),
  .y(v351)
);
assign v197 = v351;
assign v352 = v198[15:0];
assign v353 = v198[31:0];
assign v354 = v198[47:0];
assign v355 = v352[3:0];
assign v356 = (v355 == v162);
assign v357 = v352[0];
assign v358 = (~v356);
assign v359 = (v358 & v357);
assign v360 = (~v357);
assign v361 = (v358 & v360);
assign v362 = v353[11:7];
assign v363 = {{1{1'b0}}, v362};
assign v364 = v353[19:15];
assign v365 = {{1{1'b0}}, v364};
assign v366 = v353[24:20];
assign v367 = {{1{1'b0}}, v366};
assign v368 = v353[31:27];
assign v369 = {{1{1'b0}}, v368};
assign v370 = v353[31:20];
assign v371 = {{52{1'b0}}, v370};
assign v372 = {{52{v370[11]}}, v370};
assign v373 = v353[31:12];
assign v374 = {{44{v373[19]}}, v373};
assign v375 = v353[31:25];
assign v376 = {{7{1'b0}}, v362};
assign v377 = (v376 << 7);
assign v378 = {{5{1'b0}}, v375};
assign v379 = (v377 | v378);
assign v380 = {{52{v379[11]}}, v379};
assign v381 = v353[31:15];
assign v382 = {{47{v381[16]}}, v381};
assign v383 = v354[15:0];
assign v384 = v354[47:16];
assign v385 = v383[15:4];
assign v386 = v384[31:12];
assign v387 = {{20{1'b0}}, v385};
assign v388 = (v387 << 20);
assign v389 = {{12{1'b0}}, v386};
assign v390 = (v388 | v389);
assign v391 = {{32{v390[31]}}, v390};
assign v392 = v384[11:7];
assign v393 = {{1{1'b0}}, v392};
assign v394 = v352[15:11];
assign v395 = {{1{1'b0}}, v394};
assign v396 = v352[10:6];
assign v397 = {{1{1'b0}}, v396};
assign v398 = {{59{v394[4]}}, v394};
assign v399 = {{59{v396[4]}}, v396};
assign v400 = v352[15:4];
assign v401 = {{52{v400[11]}}, v400};
assign v402 = {{59{1'b0}}, v396};
assign v403 = v352[13:11];
assign v404 = {{61{1'b0}}, v403};
assign v405 = (v352 & v161);
assign v406 = (v405 == v160);
assign v407 = (v361 & v406);
assign v408 = (v407 ? v159 : v175);
assign v409 = (v407 ? v168 : v174);
assign v410 = (v407 ? v395 : v170);
assign v411 = (v407 ? v170 : v170);
assign v412 = (v407 ? v399 : v177);
assign v413 = (v352 & v158);
assign v414 = (v413 == v157);
assign v415 = (v361 & v414);
assign v416 = (v402 << 1);
assign v417 = (v415 ? v155 : v408);
assign v418 = (v415 ? v168 : v409);
assign v419 = (v415 ? v156 : v410);
assign v420 = (v415 ? v170 : v411);
assign v421 = (v415 ? v416 : v412);
assign v422 = (v405 == v154);
assign v423 = (v361 & v422);
assign v424 = (v423 ? v152 : v417);
assign v425 = (v423 ? v168 : v418);
assign v426 = (v423 ? v170 : v419);
assign v427 = (v423 ? v397 : v420);
assign v428 = (v423 ? v153 : v420);
assign v429 = (v423 ? v170 : v420);
assign v430 = (v423 ? v398 : v421);
assign v431 = (v405 == v151);
assign v432 = (v361 & v431);
assign v433 = (v432 ? v150 : v424);
assign v434 = (v432 ? v168 : v425);
assign v435 = (v432 ? v170 : v426);
assign v436 = (v432 ? v397 : v427);
assign v437 = (v432 ? v170 : v428);
assign v438 = (v432 ? v170 : v429);
assign v439 = (v432 ? v398 : v430);
assign v440 = (v405 == v149);
assign v441 = (v361 & v440);
assign v442 = (v441 ? v148 : v433);
assign v443 = (v441 ? v168 : v434);
assign v444 = (v441 ? v395 : v435);
assign v445 = (v441 ? v397 : v436);
assign v446 = (v441 ? v170 : v437);
assign v447 = (v441 ? v170 : v438);
assign v448 = (v441 ? v177 : v439);
assign v449 = (v405 == v147);
assign v450 = (v361 & v449);
assign v451 = (v450 ? v146 : v442);
assign v452 = (v450 ? v168 : v443);
assign v453 = (v450 ? v170 : v444);
assign v454 = (v450 ? v397 : v445);
assign v455 = (v450 ? v395 : v446);
assign v456 = (v450 ? v170 : v447);
assign v457 = (v450 ? v177 : v448);
assign v458 = (v413 == v145);
assign v459 = (v361 & v458);
assign v460 = (v459 ? v153 : v451);
assign v461 = (v459 ? v168 : v452);
assign v462 = (v459 ? v170 : v453);
assign v463 = (v459 ? v397 : v454);
assign v464 = (v459 ? v170 : v455);
assign v465 = (v459 ? v170 : v456);
assign v466 = (v459 ? v177 : v457);
assign v467 = (v352 & v144);
assign v468 = (v467 == v143);
assign v469 = (v361 & v468);
assign v470 = (v401 << 1);
assign v471 = (v469 ? v142 : v460);
assign v472 = (v469 ? v168 : v461);
assign v473 = (v469 ? v170 : v462);
assign v474 = (v469 ? v170 : v463);
assign v475 = (v469 ? v170 : v464);
assign v476 = (v469 ? v170 : v465);
assign v477 = (v469 ? v470 : v466);
assign v478 = (v352 & v141);
assign v479 = (v478 == v140);
assign v480 = (v361 & v479);
assign v481 = (v480 ? v139 : v471);
assign v482 = (v480 ? v168 : v472);
assign v483 = (v480 ? v170 : v473);
assign v484 = (v480 ? v170 : v474);
assign v485 = (v480 ? v170 : v475);
assign v486 = (v480 ? v170 : v476);
assign v487 = (v480 ? v404 : v477);
assign v488 = (v352 & v138);
assign v489 = (v488 == v140);
assign v490 = (v361 & v489);
assign v491 = (v490 ? v137 : v481);
assign v492 = (v490 ? v168 : v482);
assign v493 = (v490 ? v170 : v483);
assign v494 = (v490 ? v170 : v484);
assign v495 = (v490 ? v170 : v485);
assign v496 = (v490 ? v170 : v486);
assign v497 = (v490 ? v177 : v487);
assign v498 = (v353 & v136);
assign v499 = (v498 == v135);
assign v500 = (v359 & v499);
assign v501 = (v500 ? v134 : v491);
assign v502 = (v500 ? v166 : v492);
assign v503 = (v500 ? v363 : v493);
assign v504 = (v500 ? v365 : v494);
assign v505 = (v500 ? v367 : v495);
assign v506 = (v500 ? v170 : v496);
assign v507 = (v500 ? v177 : v497);
assign v508 = (v498 == v133);
assign v509 = (v359 & v508);
assign v510 = (v509 ? v132 : v501);
assign v511 = (v509 ? v166 : v502);
assign v512 = (v509 ? v363 : v503);
assign v513 = (v509 ? v365 : v504);
assign v514 = (v509 ? v367 : v505);
assign v515 = (v509 ? v170 : v506);
assign v516 = (v509 ? v177 : v507);
assign v517 = (v498 == v131);
assign v518 = (v359 & v517);
assign v519 = (v518 ? v130 : v510);
assign v520 = (v518 ? v166 : v511);
assign v521 = (v518 ? v363 : v512);
assign v522 = (v518 ? v365 : v513);
assign v523 = (v518 ? v367 : v514);
assign v524 = (v518 ? v170 : v515);
assign v525 = (v518 ? v177 : v516);
assign v526 = (v498 == v129);
assign v527 = (v359 & v526);
assign v528 = (v527 ? v128 : v519);
assign v529 = (v527 ? v166 : v520);
assign v530 = (v527 ? v363 : v521);
assign v531 = (v527 ? v365 : v522);
assign v532 = (v527 ? v367 : v523);
assign v533 = (v527 ? v170 : v524);
assign v534 = (v527 ? v177 : v525);
assign v535 = (v498 == v127);
assign v536 = (v359 & v535);
assign v537 = (v536 ? v126 : v528);
assign v538 = (v536 ? v166 : v529);
assign v539 = (v536 ? v363 : v530);
assign v540 = (v536 ? v365 : v531);
assign v541 = (v536 ? v367 : v532);
assign v542 = (v536 ? v369 : v533);
assign v543 = (v536 ? v177 : v534);
assign v544 = (v498 == v125);
assign v545 = (v359 & v544);
assign v546 = (v545 ? v156 : v537);
assign v547 = (v545 ? v166 : v538);
assign v548 = (v545 ? v170 : v539);
assign v549 = (v545 ? v365 : v540);
assign v550 = (v545 ? v367 : v541);
assign v551 = (v545 ? v170 : v542);
assign v552 = (v545 ? v380 : v543);
assign v553 = (v498 == v124);
assign v554 = (v359 & v553);
assign v555 = (v554 ? v123 : v546);
assign v556 = (v554 ? v166 : v547);
assign v557 = (v554 ? v170 : v548);
assign v558 = (v554 ? v365 : v549);
assign v559 = (v554 ? v367 : v550);
assign v560 = (v554 ? v170 : v551);
assign v561 = (v554 ? v380 : v552);
assign v562 = (v498 == v122);
assign v563 = (v359 & v562);
assign v564 = (v563 ? v121 : v555);
assign v565 = (v563 ? v166 : v556);
assign v566 = (v563 ? v363 : v557);
assign v567 = (v563 ? v365 : v558);
assign v568 = (v563 ? v170 : v559);
assign v569 = (v563 ? v170 : v560);
assign v570 = (v563 ? v372 : v561);
assign v571 = (v498 == v120);
assign v572 = (v359 & v571);
assign v573 = (v572 ? v119 : v564);
assign v574 = (v572 ? v166 : v565);
assign v575 = (v572 ? v363 : v566);
assign v576 = (v572 ? v365 : v567);
assign v577 = (v572 ? v170 : v568);
assign v578 = (v572 ? v170 : v569);
assign v579 = (v572 ? v371 : v570);
assign v580 = (v498 == v118);
assign v581 = (v359 & v580);
assign v582 = (v581 ? v117 : v573);
assign v583 = (v581 ? v166 : v574);
assign v584 = (v581 ? v363 : v575);
assign v585 = (v581 ? v365 : v576);
assign v586 = (v581 ? v170 : v577);
assign v587 = (v581 ? v170 : v578);
assign v588 = (v581 ? v371 : v579);
assign v589 = (v498 == v116);
assign v590 = (v359 & v589);
assign v591 = (v590 ? v115 : v582);
assign v592 = (v590 ? v166 : v583);
assign v593 = (v590 ? v363 : v584);
assign v594 = (v590 ? v365 : v585);
assign v595 = (v590 ? v170 : v586);
assign v596 = (v590 ? v170 : v587);
assign v597 = (v590 ? v371 : v588);
assign v598 = (v353 & v114);
assign v599 = (v598 == v113);
assign v600 = (v359 & v599);
assign v601 = (v600 ? v112 : v591);
assign v602 = (v600 ? v166 : v592);
assign v603 = (v600 ? v363 : v593);
assign v604 = (v600 ? v365 : v594);
assign v605 = (v600 ? v367 : v595);
assign v606 = (v600 ? v170 : v596);
assign v607 = (v600 ? v177 : v597);
assign v608 = (v353 & v111);
assign v609 = (v608 == v110);
assign v610 = (v359 & v609);
assign v611 = (v610 ? v165 : v601);
assign v612 = (v610 ? v166 : v602);
assign v613 = (v610 ? v170 : v603);
assign v614 = (v610 ? v170 : v604);
assign v615 = (v610 ? v170 : v605);
assign v616 = (v610 ? v170 : v606);
assign v617 = (v610 ? v177 : v607);
assign v618 = (v353 & v109);
assign v619 = (v618 == v108);
assign v620 = (v359 & v619);
assign v621 = (v374 << 12);
assign v622 = (v620 ? v107 : v611);
assign v623 = (v620 ? v166 : v612);
assign v624 = (v620 ? v363 : v613);
assign v625 = (v620 ? v170 : v614);
assign v626 = (v620 ? v170 : v615);
assign v627 = (v620 ? v170 : v616);
assign v628 = (v620 ? v621 : v617);
assign v629 = (v353 & v106);
assign v630 = (v629 == v105);
assign v631 = (v359 & v630);
assign v632 = (v382 << 1);
assign v633 = (v631 ? v104 : v622);
assign v634 = (v631 ? v166 : v623);
assign v635 = (v631 ? v170 : v624);
assign v636 = (v631 ? v170 : v625);
assign v637 = (v631 ? v170 : v626);
assign v638 = (v631 ? v170 : v627);
assign v639 = (v631 ? v632 : v628);
assign v640 = (v354 & v103);
assign v641 = (v640 == v102);
assign v642 = (v356 & v641);
assign v643 = (v642 ? v101 : v633);
assign v644 = (v642 ? v100 : v634);
assign v645 = (v642 ? v393 : v635);
assign v646 = (v642 ? v170 : v636);
assign v647 = (v642 ? v170 : v637);
assign v648 = (v642 ? v170 : v638);
assign v649 = (v642 ? v391 : v639);
assign v650 = (v343 ? v643 : v200);
assign v651 = v644;
assign v652 = v645;
assign v653 = v646;
assign v654 = v647;
assign v655 = v648;
assign v656 = v649;
assign v657 = v650;
assign v199 = v657;
pyc_mux #(.WIDTH(3)) v658_inst (
  .sel(v343),
  .a(v651),
  .b(v202),
  .y(v658)
);
assign v201 = v658;
pyc_mux #(.WIDTH(6)) v659_inst (
  .sel(v343),
  .a(v652),
  .b(v204),
  .y(v659)
);
assign v203 = v659;
pyc_mux #(.WIDTH(6)) v660_inst (
  .sel(v343),
  .a(v653),
  .b(v206),
  .y(v660)
);
assign v205 = v660;
pyc_mux #(.WIDTH(6)) v661_inst (
  .sel(v343),
  .a(v654),
  .b(v208),
  .y(v661)
);
assign v207 = v661;
pyc_mux #(.WIDTH(6)) v662_inst (
  .sel(v343),
  .a(v655),
  .b(v210),
  .y(v662)
);
assign v209 = v662;
pyc_mux #(.WIDTH(64)) v663_inst (
  .sel(v343),
  .a(v656),
  .b(v212),
  .y(v663)
);
assign v211 = v663;
assign v664 = (v653 == v175);
assign v665 = (v664 ? v177 : v177);
assign v666 = (v653 == v139);
assign v667 = (v666 ? v248 : v665);
assign v668 = (v653 == v137);
assign v669 = (v668 ? v250 : v667);
assign v670 = (v653 == v148);
assign v671 = (v670 ? v252 : v669);
assign v672 = (v653 == v150);
assign v673 = (v672 ? v254 : v671);
assign v674 = (v653 == v152);
assign v675 = (v674 ? v256 : v673);
assign v676 = (v653 == v115);
assign v677 = (v676 ? v258 : v675);
assign v678 = (v653 == v117);
assign v679 = (v678 ? v260 : v677);
assign v680 = (v653 == v119);
assign v681 = (v680 ? v262 : v679);
assign v682 = (v653 == v121);
assign v683 = (v682 ? v264 : v681);
assign v684 = (v653 == v156);
assign v685 = (v684 ? v266 : v683);
assign v686 = (v653 == v128);
assign v687 = (v686 ? v268 : v685);
assign v688 = (v653 == v130);
assign v689 = (v688 ? v270 : v687);
assign v690 = (v653 == v132);
assign v691 = (v690 ? v272 : v689);
assign v692 = (v653 == v134);
assign v693 = (v692 ? v274 : v691);
assign v694 = (v653 == v112);
assign v695 = (v694 ? v276 : v693);
assign v696 = (v653 == v126);
assign v697 = (v696 ? v278 : v695);
assign v698 = (v653 == v101);
assign v699 = (v698 ? v280 : v697);
assign v700 = (v653 == v165);
assign v701 = (v700 ? v282 : v699);
assign v702 = (v653 == v142);
assign v703 = (v702 ? v284 : v701);
assign v704 = (v653 == v104);
assign v705 = (v704 ? v286 : v703);
assign v706 = (v653 == v159);
assign v707 = (v706 ? v288 : v705);
assign v708 = (v653 == v155);
assign v709 = (v708 ? v290 : v707);
assign v710 = (v653 == v146);
assign v711 = (v710 ? v292 : v709);
assign v712 = (v653 == v153);
assign v713 = (v712 ? v294 : v711);
assign v714 = (v653 == v107);
assign v715 = (v714 ? v296 : v713);
assign v716 = (v653 == v123);
assign v717 = (v716 ? v298 : v715);
assign v718 = (v653 == v99);
assign v719 = (v718 ? v300 : v717);
assign v720 = (v653 == v98);
assign v721 = (v720 ? v302 : v719);
assign v722 = (v653 == v97);
assign v723 = (v722 ? v304 : v721);
assign v724 = (v653 == v96);
assign v725 = (v724 ? v306 : v723);
assign v726 = (v653 == v95);
assign v727 = (v726 ? v308 : v725);
assign v728 = (v654 == v175);
assign v729 = (v728 ? v177 : v177);
assign v730 = (v654 == v139);
assign v731 = (v730 ? v248 : v729);
assign v732 = (v654 == v137);
assign v733 = (v732 ? v250 : v731);
assign v734 = (v654 == v148);
assign v735 = (v734 ? v252 : v733);
assign v736 = (v654 == v150);
assign v737 = (v736 ? v254 : v735);
assign v738 = (v654 == v152);
assign v739 = (v738 ? v256 : v737);
assign v740 = (v654 == v115);
assign v741 = (v740 ? v258 : v739);
assign v742 = (v654 == v117);
assign v743 = (v742 ? v260 : v741);
assign v744 = (v654 == v119);
assign v745 = (v744 ? v262 : v743);
assign v746 = (v654 == v121);
assign v747 = (v746 ? v264 : v745);
assign v748 = (v654 == v156);
assign v749 = (v748 ? v266 : v747);
assign v750 = (v654 == v128);
assign v751 = (v750 ? v268 : v749);
assign v752 = (v654 == v130);
assign v753 = (v752 ? v270 : v751);
assign v754 = (v654 == v132);
assign v755 = (v754 ? v272 : v753);
assign v756 = (v654 == v134);
assign v757 = (v756 ? v274 : v755);
assign v758 = (v654 == v112);
assign v759 = (v758 ? v276 : v757);
assign v760 = (v654 == v126);
assign v761 = (v760 ? v278 : v759);
assign v762 = (v654 == v101);
assign v763 = (v762 ? v280 : v761);
assign v764 = (v654 == v165);
assign v765 = (v764 ? v282 : v763);
assign v766 = (v654 == v142);
assign v767 = (v766 ? v284 : v765);
assign v768 = (v654 == v104);
assign v769 = (v768 ? v286 : v767);
assign v770 = (v654 == v159);
assign v771 = (v770 ? v288 : v769);
assign v772 = (v654 == v155);
assign v773 = (v772 ? v290 : v771);
assign v774 = (v654 == v146);
assign v775 = (v774 ? v292 : v773);
assign v776 = (v654 == v153);
assign v777 = (v776 ? v294 : v775);
assign v778 = (v654 == v107);
assign v779 = (v778 ? v296 : v777);
assign v780 = (v654 == v123);
assign v781 = (v780 ? v298 : v779);
assign v782 = (v654 == v99);
assign v783 = (v782 ? v300 : v781);
assign v784 = (v654 == v98);
assign v785 = (v784 ? v302 : v783);
assign v786 = (v654 == v97);
assign v787 = (v786 ? v304 : v785);
assign v788 = (v654 == v96);
assign v789 = (v788 ? v306 : v787);
assign v790 = (v654 == v95);
assign v791 = (v790 ? v308 : v789);
assign v792 = (v655 == v175);
assign v793 = (v792 ? v177 : v177);
assign v794 = (v655 == v139);
assign v795 = (v794 ? v248 : v793);
assign v796 = (v655 == v137);
assign v797 = (v796 ? v250 : v795);
assign v798 = (v655 == v148);
assign v799 = (v798 ? v252 : v797);
assign v800 = (v655 == v150);
assign v801 = (v800 ? v254 : v799);
assign v802 = (v655 == v152);
assign v803 = (v802 ? v256 : v801);
assign v804 = (v655 == v115);
assign v805 = (v804 ? v258 : v803);
assign v806 = (v655 == v117);
assign v807 = (v806 ? v260 : v805);
assign v808 = (v655 == v119);
assign v809 = (v808 ? v262 : v807);
assign v810 = (v655 == v121);
assign v811 = (v810 ? v264 : v809);
assign v812 = (v655 == v156);
assign v813 = (v812 ? v266 : v811);
assign v814 = (v655 == v128);
assign v815 = (v814 ? v268 : v813);
assign v816 = (v655 == v130);
assign v817 = (v816 ? v270 : v815);
assign v818 = (v655 == v132);
assign v819 = (v818 ? v272 : v817);
assign v820 = (v655 == v134);
assign v821 = (v820 ? v274 : v819);
assign v822 = (v655 == v112);
assign v823 = (v822 ? v276 : v821);
assign v824 = (v655 == v126);
assign v825 = (v824 ? v278 : v823);
assign v826 = (v655 == v101);
assign v827 = (v826 ? v280 : v825);
assign v828 = (v655 == v165);
assign v829 = (v828 ? v282 : v827);
assign v830 = (v655 == v142);
assign v831 = (v830 ? v284 : v829);
assign v832 = (v655 == v104);
assign v833 = (v832 ? v286 : v831);
assign v834 = (v655 == v159);
assign v835 = (v834 ? v288 : v833);
assign v836 = (v655 == v155);
assign v837 = (v836 ? v290 : v835);
assign v838 = (v655 == v146);
assign v839 = (v838 ? v292 : v837);
assign v840 = (v655 == v153);
assign v841 = (v840 ? v294 : v839);
assign v842 = (v655 == v107);
assign v843 = (v842 ? v296 : v841);
assign v844 = (v655 == v123);
assign v845 = (v844 ? v298 : v843);
assign v846 = (v655 == v99);
assign v847 = (v846 ? v300 : v845);
assign v848 = (v655 == v98);
assign v849 = (v848 ? v302 : v847);
assign v850 = (v655 == v97);
assign v851 = (v850 ? v304 : v849);
assign v852 = (v655 == v96);
assign v853 = (v852 ? v306 : v851);
assign v854 = (v655 == v95);
assign v855 = (v854 ? v308 : v853);
assign v856 = (v343 ? v727 : v214);
assign v857 = v791;
assign v858 = v855;
assign v859 = v856;
assign v213 = v859;
pyc_mux #(.WIDTH(64)) v860_inst (
  .sel(v343),
  .a(v857),
  .b(v216),
  .y(v860)
);
assign v215 = v860;
pyc_mux #(.WIDTH(64)) v861_inst (
  .sel(v343),
  .a(v858),
  .b(v218),
  .y(v861)
);
assign v217 = v861;
assign v862 = (v200 == v139);
assign v863 = (v200 == v142);
assign v864 = (v200 == v104);
assign v865 = (v200 == v148);
assign v866 = (v200 == v159);
assign v867 = (v200 == v155);
assign v868 = (v200 == v146);
assign v869 = (v200 == v153);
assign v870 = (v200 == v107);
assign v871 = (v200 == v117);
assign v872 = (v200 == v115);
assign v873 = (v200 == v119);
assign v874 = (v200 == v128);
assign v875 = (v200 == v130);
assign v876 = (v200 == v132);
assign v877 = (v200 == v134);
assign v878 = (v200 == v112);
assign v879 = (v200 == v126);
assign v880 = (v200 == v101);
assign v881 = (v200 == v121);
assign v882 = (v200 == v150);
assign v883 = (v200 == v156);
assign v884 = (v200 == v152);
assign v885 = (v200 == v123);
assign v886 = (v212 << 2);
assign v887 = (v862 | v863);
assign v888 = (v887 | v864);
assign v889 = (v888 ? v212 : v177);
assign v890 = (v888 ? v173 : v173);
assign v891 = (v888 ? v174 : v174);
assign v892 = (v888 ? v177 : v177);
assign v893 = (v865 ? v214 : v889);
assign v894 = (v865 ? v173 : v890);
assign v895 = (v865 ? v174 : v891);
assign v896 = (v865 ? v177 : v892);
assign v897 = (v866 ? v212 : v893);
assign v898 = (v866 ? v173 : v894);
assign v899 = (v866 ? v174 : v895);
assign v900 = (v866 ? v177 : v896);
assign v901 = (v182 + v212);
assign v902 = (v867 ? v901 : v897);
assign v903 = (v867 ? v173 : v898);
assign v904 = (v867 ? v174 : v899);
assign v905 = (v867 ? v177 : v900);
assign v906 = (v214 == v216);
assign v907 = (v906 ? v178 : v177);
assign v908 = (v868 ? v907 : v902);
assign v909 = (v868 ? v173 : v903);
assign v910 = (v868 ? v174 : v904);
assign v911 = (v868 ? v177 : v905);
assign v912 = (v869 ? v214 : v908);
assign v913 = (v869 ? v173 : v909);
assign v914 = (v869 ? v174 : v910);
assign v915 = (v869 ? v177 : v911);
assign v916 = (v182 & v94);
assign v917 = (v916 + v212);
assign v918 = (v870 ? v917 : v912);
assign v919 = (v870 ? v173 : v913);
assign v920 = (v870 ? v174 : v914);
assign v921 = (v870 ? v177 : v915);
assign v922 = (v214 + v212);
assign v923 = (v871 ? v922 : v918);
assign v924 = (v871 ? v173 : v919);
assign v925 = (v871 ? v174 : v920);
assign v926 = (v871 ? v177 : v921);
assign v927 = (~v212);
assign v928 = (v927 + v178);
assign v929 = (v214 + v928);
assign v930 = (v872 ? v929 : v923);
assign v931 = (v872 ? v173 : v924);
assign v932 = (v872 ? v174 : v925);
assign v933 = (v872 ? v177 : v926);
assign v934 = v214[31:0];
assign v935 = v212[31:0];
assign v936 = (v934 + v935);
assign v937 = {{32{v936[31]}}, v936};
assign v938 = (v873 ? v937 : v930);
assign v939 = (v873 ? v173 : v931);
assign v940 = (v873 ? v174 : v932);
assign v941 = (v873 ? v177 : v933);
assign v942 = v216[31:0];
assign v943 = (v934 + v942);
assign v944 = {{32{v943[31]}}, v943};
assign v945 = (v934 | v942);
assign v946 = {{32{v945[31]}}, v945};
assign v947 = (v934 & v942);
assign v948 = {{32{v947[31]}}, v947};
assign v949 = (v934 ^ v942);
assign v950 = {{32{v949[31]}}, v949};
assign v951 = (v874 ? v944 : v938);
assign v952 = (v874 ? v173 : v939);
assign v953 = (v874 ? v174 : v940);
assign v954 = (v874 ? v177 : v941);
assign v955 = (v875 ? v946 : v951);
assign v956 = (v875 ? v173 : v952);
assign v957 = (v875 ? v174 : v953);
assign v958 = (v875 ? v177 : v954);
assign v959 = (v876 ? v948 : v955);
assign v960 = (v876 ? v173 : v956);
assign v961 = (v876 ? v174 : v957);
assign v962 = (v876 ? v177 : v958);
assign v963 = (v877 ? v950 : v959);
assign v964 = (v877 ? v173 : v960);
assign v965 = (v877 ? v174 : v961);
assign v966 = (v877 ? v177 : v962);
assign v967 = (v878 ? v907 : v963);
assign v968 = (v878 ? v173 : v964);
assign v969 = (v878 ? v174 : v965);
assign v970 = (v878 ? v177 : v966);
assign v971 = (v880 ? v212 : v967);
assign v972 = (v880 ? v173 : v968);
assign v973 = (v880 ? v174 : v969);
assign v974 = (v880 ? v177 : v970);
assign v975 = (v218 == v177);
assign v976 = (~v975);
assign v977 = (v976 ? v216 : v214);
assign v978 = (v879 ? v977 : v971);
assign v979 = (v879 ? v173 : v972);
assign v980 = (v879 ? v174 : v973);
assign v981 = (v879 ? v177 : v974);
assign v982 = (v881 | v882);
assign v983 = (v214 + v886);
assign v984 = (v982 ? v177 : v978);
assign v985 = (v982 ? v172 : v979);
assign v986 = (v982 ? v173 : v979);
assign v987 = (v982 ? v166 : v980);
assign v988 = (v982 ? v983 : v981);
assign v989 = (v982 ? v177 : v981);
assign v990 = (v216 + v886);
assign v991 = (v883 ? v990 : v983);
assign v992 = (v883 ? v214 : v216);
assign v993 = (v883 | v884);
assign v994 = (v993 ? v177 : v984);
assign v995 = (v993 ? v173 : v985);
assign v996 = (v993 ? v172 : v986);
assign v997 = (v993 ? v166 : v987);
assign v998 = (v993 ? v991 : v988);
assign v999 = (v993 ? v992 : v989);
assign v1000 = (v212 << 3);
assign v1001 = (v216 + v1000);
assign v1002 = (v885 ? v177 : v994);
assign v1003 = (v885 ? v173 : v995);
assign v1004 = (v885 ? v172 : v996);
assign v1005 = (v885 ? v174 : v997);
assign v1006 = (v885 ? v1001 : v998);
assign v1007 = (v885 ? v214 : v999);
assign v1008 = (v344 ? v200 : v220);
assign v1009 = v1002;
assign v1010 = v1003;
assign v1011 = v1004;
assign v1012 = v1005;
assign v1013 = v1006;
assign v1014 = v1007;
assign v1015 = v1008;
assign v219 = v1015;
pyc_mux #(.WIDTH(3)) v1016_inst (
  .sel(v344),
  .a(v202),
  .b(v222),
  .y(v1016)
);
assign v221 = v1016;
pyc_mux #(.WIDTH(6)) v1017_inst (
  .sel(v344),
  .a(v204),
  .b(v224),
  .y(v1017)
);
assign v223 = v1017;
pyc_mux #(.WIDTH(64)) v1018_inst (
  .sel(v344),
  .a(v1009),
  .b(v226),
  .y(v1018)
);
assign v225 = v1018;
pyc_mux #(.WIDTH(1)) v1019_inst (
  .sel(v344),
  .a(v1010),
  .b(v228),
  .y(v1019)
);
assign v227 = v1019;
pyc_mux #(.WIDTH(1)) v1020_inst (
  .sel(v344),
  .a(v1011),
  .b(v230),
  .y(v1020)
);
assign v229 = v1020;
pyc_mux #(.WIDTH(3)) v1021_inst (
  .sel(v344),
  .a(v1012),
  .b(v232),
  .y(v1021)
);
assign v231 = v1021;
pyc_mux #(.WIDTH(64)) v1022_inst (
  .sel(v344),
  .a(v1013),
  .b(v234),
  .y(v1022)
);
assign v233 = v1022;
pyc_mux #(.WIDTH(64)) v1023_inst (
  .sel(v344),
  .a(v1014),
  .b(v236),
  .y(v1023)
);
assign v235 = v1023;
assign v1024 = v350[31:0];
assign v1025 = {{32{v1024[31]}}, v1024};
assign v1026 = (v228 ? v1025 : v226);
assign v1027 = (v230 ? v177 : v1026);
assign v1028 = (v345 ? v220 : v238);
assign v1029 = v1027;
assign v1030 = v1028;
assign v237 = v1030;
pyc_mux #(.WIDTH(3)) v1031_inst (
  .sel(v345),
  .a(v222),
  .b(v240),
  .y(v1031)
);
assign v239 = v1031;
pyc_mux #(.WIDTH(6)) v1032_inst (
  .sel(v345),
  .a(v224),
  .b(v242),
  .y(v1032)
);
assign v241 = v1032;
pyc_mux #(.WIDTH(64)) v1033_inst (
  .sel(v345),
  .a(v1029),
  .b(v244),
  .y(v1033)
);
assign v243 = v1033;
pyc_mux #(.WIDTH(1)) v1034_inst (
  .sel(v340),
  .a(v172),
  .b(v196),
  .y(v1034)
);
assign v195 = v1034;
assign v1035 = (v238 == v139);
assign v1036 = (v238 == v142);
assign v1037 = (v238 == v104);
assign v1038 = (v238 == v137);
assign v1039 = (v1035 | v1036);
assign v1040 = (v1039 | v1037);
assign v1041 = (v1040 | v1038);
assign v1042 = (v184 == v93);
assign v1043 = (v184 == v92);
assign v1044 = (v184 == v91);
assign v1045 = (v186 + v188);
assign v1046 = (v1044 ? v192 : v1045);
assign v1047 = (v1043 | v1044);
assign v1048 = (v1042 & v190);
assign v1049 = (v1047 | v1048);
assign v1050 = {{61{1'b0}}, v240};
assign v1051 = (v182 + v1050);
assign v1052 = (v1049 ? v1046 : v1051);
assign v1053 = (v1041 ? v1052 : v1051);
assign v1054 = (v346 ? v1053 : v182);
assign v1055 = v1035;
assign v1056 = v1036;
assign v1057 = v1037;
assign v1058 = v1038;
assign v1059 = v1040;
assign v1060 = v1041;
assign v1061 = v1049;
assign v1062 = v1054;
assign v181 = v1062;
assign v1063 = (v335 ? v169 : v180);
assign v1064 = (v336 ? v168 : v1063);
assign v1065 = (v337 ? v167 : v1064);
assign v1066 = (v338 ? v166 : v1065);
assign v1067 = (v339 ? v174 : v1066);
assign v1068 = (v341 ? v180 : v1067);
assign v1069 = v1068;
assign v179 = v1069;
pyc_add #(.WIDTH(64)) v1070_inst (
  .a(v194),
  .b(v178),
  .y(v1070)
);
assign v193 = v1070;
assign v1071 = (v238 == v146);
assign v1072 = (v238 == v153);
assign v1073 = (v346 & v1060);
assign v1074 = (v1073 ? v173 : v190);
assign v1075 = (v1073 ? v177 : v192);
assign v1076 = (v346 & v1071);
assign v1077 = v244[0];
assign v1078 = (v1076 ? v1077 : v1074);
assign v1079 = (v346 & v1072);
assign v1080 = (v1079 ? v244 : v1075);
assign v1081 = v1073;
assign v1082 = v1078;
assign v1083 = v1080;
assign v189 = v1082;
assign v191 = v1083;
assign v1084 = (v1081 & v1061);
assign v1085 = (v1084 ? v171 : v184);
assign v1086 = (v1084 ? v182 : v186);
assign v1087 = (v1084 ? v177 : v188);
assign v1088 = (v346 & v1059);
assign v1089 = (~v1061);
assign v1090 = (v1088 & v1089);
assign v1091 = (v1090 & v1056);
assign v1092 = (v1091 ? v93 : v1085);
assign v1093 = (v1091 ? v182 : v1086);
assign v1094 = (v1091 ? v244 : v1087);
assign v1095 = (v1090 & v1057);
assign v1096 = (v1095 ? v92 : v1092);
assign v1097 = (v1095 ? v182 : v1093);
assign v1098 = (v1095 ? v244 : v1094);
assign v1099 = v244[2:0];
assign v1100 = (v1099 == v90);
assign v1101 = (v1100 ? v91 : v171);
assign v1102 = (v1090 & v1055);
assign v1103 = (v1102 ? v1101 : v1096);
assign v1104 = (v1102 ? v182 : v1097);
assign v1105 = (v1102 ? v177 : v1098);
assign v1106 = (v346 & v1058);
assign v1107 = (v1106 ? v171 : v1103);
assign v1108 = (v1106 ? v182 : v1104);
assign v1109 = (v1106 ? v177 : v1105);
assign v1110 = v1088;
assign v1111 = v1107;
assign v1112 = v1108;
assign v1113 = v1109;
assign v183 = v1111;
assign v185 = v1112;
assign v187 = v1113;
assign v1114 = (v238 == v156);
assign v1115 = (v238 == v152);
assign v1116 = (v1114 | v1115);
assign v1117 = (~v1116);
assign v1118 = (v346 & v1117);
assign v1119 = (v242 == v170);
assign v1120 = (~v1119);
assign v1121 = (v1118 & v1120);
assign v1122 = (v238 == v150);
assign v1123 = (v346 & v1122);
assign v1124 = (v242 == v95);
assign v1125 = (v1121 & v1124);
assign v1126 = (v1123 | v1125);
assign v1127 = (v242 == v96);
assign v1128 = (v1121 & v1127);
assign v1129 = v1121;
assign v1130 = v1126;
assign v1131 = v1128;
assign v245 = v177;
assign v1132 = (v242 == v139);
assign v1133 = (v1129 & v1132);
assign v1134 = (v1133 ? v244 : v248);
assign v1135 = v1134;
assign v247 = v1135;
assign v1136 = (v242 == v137);
assign v1137 = (v1129 & v1136);
assign v1138 = (v1137 ? v244 : v250);
assign v1139 = v1138;
assign v249 = v1139;
assign v1140 = (v242 == v148);
assign v1141 = (v1129 & v1140);
assign v1142 = (v1141 ? v244 : v252);
assign v1143 = v1142;
assign v251 = v1143;
assign v1144 = (v242 == v150);
assign v1145 = (v1129 & v1144);
assign v1146 = (v1145 ? v244 : v254);
assign v1147 = v1146;
assign v253 = v1147;
assign v1148 = (v242 == v152);
assign v1149 = (v1129 & v1148);
assign v1150 = (v1149 ? v244 : v256);
assign v1151 = v1150;
assign v255 = v1151;
assign v1152 = (v242 == v115);
assign v1153 = (v1129 & v1152);
assign v1154 = (v1153 ? v244 : v258);
assign v1155 = v1154;
assign v257 = v1155;
assign v1156 = (v242 == v117);
assign v1157 = (v1129 & v1156);
assign v1158 = (v1157 ? v244 : v260);
assign v1159 = v1158;
assign v259 = v1159;
assign v1160 = (v242 == v119);
assign v1161 = (v1129 & v1160);
assign v1162 = (v1161 ? v244 : v262);
assign v1163 = v1162;
assign v261 = v1163;
assign v1164 = (v242 == v121);
assign v1165 = (v1129 & v1164);
assign v1166 = (v1165 ? v244 : v264);
assign v1167 = v1166;
assign v263 = v1167;
assign v1168 = (v242 == v156);
assign v1169 = (v1129 & v1168);
assign v1170 = (v1169 ? v244 : v266);
assign v1171 = v1170;
assign v265 = v1171;
assign v1172 = (v242 == v128);
assign v1173 = (v1129 & v1172);
assign v1174 = (v1173 ? v244 : v268);
assign v1175 = v1174;
assign v267 = v1175;
assign v1176 = (v242 == v130);
assign v1177 = (v1129 & v1176);
assign v1178 = (v1177 ? v244 : v270);
assign v1179 = v1178;
assign v269 = v1179;
assign v1180 = (v242 == v132);
assign v1181 = (v1129 & v1180);
assign v1182 = (v1181 ? v244 : v272);
assign v1183 = v1182;
assign v271 = v1183;
assign v1184 = (v242 == v134);
assign v1185 = (v1129 & v1184);
assign v1186 = (v1185 ? v244 : v274);
assign v1187 = v1186;
assign v273 = v1187;
assign v1188 = (v242 == v112);
assign v1189 = (v1129 & v1188);
assign v1190 = (v1189 ? v244 : v276);
assign v1191 = v1190;
assign v275 = v1191;
assign v1192 = (v242 == v126);
assign v1193 = (v1129 & v1192);
assign v1194 = (v1193 ? v244 : v278);
assign v1195 = v1194;
assign v277 = v1195;
assign v1196 = (v242 == v101);
assign v1197 = (v1129 & v1196);
assign v1198 = (v1197 ? v244 : v280);
assign v1199 = v1198;
assign v279 = v1199;
assign v1200 = (v242 == v165);
assign v1201 = (v1129 & v1200);
assign v1202 = (v1201 ? v244 : v282);
assign v1203 = v1202;
assign v281 = v1203;
assign v1204 = (v242 == v142);
assign v1205 = (v1129 & v1204);
assign v1206 = (v1205 ? v244 : v284);
assign v1207 = v1206;
assign v283 = v1207;
assign v1208 = (v242 == v104);
assign v1209 = (v1129 & v1208);
assign v1210 = (v1209 ? v244 : v286);
assign v1211 = v1210;
assign v285 = v1211;
assign v1212 = (v242 == v159);
assign v1213 = (v1129 & v1212);
assign v1214 = (v1213 ? v244 : v288);
assign v1215 = v1214;
assign v287 = v1215;
assign v1216 = (v242 == v155);
assign v1217 = (v1129 & v1216);
assign v1218 = (v1217 ? v244 : v290);
assign v1219 = v1218;
assign v289 = v1219;
assign v1220 = (v242 == v146);
assign v1221 = (v1129 & v1220);
assign v1222 = (v1221 ? v244 : v292);
assign v1223 = v1222;
assign v291 = v1223;
assign v1224 = (v1130 ? v244 : v294);
assign v1225 = (v1110 ? v177 : v1224);
assign v1226 = (v1130 ? v294 : v296);
assign v1227 = (v1110 ? v177 : v1226);
assign v1228 = (v1130 ? v296 : v298);
assign v1229 = (v1110 ? v177 : v1228);
assign v1230 = (v1130 ? v298 : v300);
assign v1231 = (v1110 ? v177 : v1230);
assign v1232 = (v1131 ? v244 : v302);
assign v1233 = (v1110 ? v177 : v1232);
assign v1234 = (v1131 ? v302 : v304);
assign v1235 = (v1110 ? v177 : v1234);
assign v1236 = (v1131 ? v304 : v306);
assign v1237 = (v1110 ? v177 : v1236);
assign v1238 = (v1131 ? v306 : v308);
assign v1239 = (v1110 ? v177 : v1238);
assign v1240 = v1225;
assign v1241 = v1227;
assign v1242 = v1229;
assign v1243 = v1231;
assign v1244 = v1233;
assign v1245 = v1235;
assign v1246 = v1237;
assign v1247 = v1239;
assign v293 = v1240;
assign v295 = v1241;
assign v297 = v1242;
assign v299 = v1243;
assign v301 = v1244;
assign v303 = v1245;
assign v305 = v1246;
assign v307 = v1247;
assign halted = v196;
assign pc = v182;
assign stage = v180;
assign cycles = v194;
assign a0 = v250;
assign a1 = v252;
assign ra = v266;
assign sp = v248;
assign br_kind = v184;
assign if_window = v198;
assign wb_op = v238;
assign wb_regdst = v242;
assign wb_value = v244;
assign commit_cond = v190;
assign commit_tgt = v192;

endmodule

